module Nand(
	input a,
	input b,
	output out
);

	nand(out, a, b);

endmodule
